module notGate(a, inversedA);

input a;
output inversedA;

assign inversedA = ~a;

endmodule