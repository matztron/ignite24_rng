module inv (
    input i,
    output q
);

assign q = ~i;

endmodule